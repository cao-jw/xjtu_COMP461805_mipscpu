module Add1(
    A,B,C
    );
    input [31:0] A,B;
    output [31:0] C;
    assign C = A + B;
endmodule
