module OrGate(A,B,R);
input A,B;
output R;
assign R=A|B;
endmodule