module AndGate(
R,A,B
    );
    input A,B;
    output  R;
    assign R=A&B;
endmodule
